VERSION 5.4 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
  DATABASE MICRONS 2000 ;
END UNITS
MACRO sram_32b_256_1rw_sky130
   CLASS BLOCK ;
   SIZE 288.94 BY 502.86 ;
   SYMMETRY X Y R90 ;
   PIN din0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  78.8 0.0 79.18 0.38 ;
      END
   END din0[0]
   PIN din0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  84.64 0.0 85.02 0.38 ;
      END
   END din0[1]
   PIN din0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  90.48 0.0 90.86 0.38 ;
      END
   END din0[2]
   PIN din0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  96.32 0.0 96.7 0.38 ;
      END
   END din0[3]
   PIN din0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  102.16 0.0 102.54 0.38 ;
      END
   END din0[4]
   PIN din0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  108.0 0.0 108.38 0.38 ;
      END
   END din0[5]
   PIN din0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  113.84 0.0 114.22 0.38 ;
      END
   END din0[6]
   PIN din0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  119.68 0.0 120.06 0.38 ;
      END
   END din0[7]
   PIN din0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  125.52 0.0 125.9 0.38 ;
      END
   END din0[8]
   PIN din0[9]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  131.36 0.0 131.74 0.38 ;
      END
   END din0[9]
   PIN din0[10]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  137.2 0.0 137.58 0.38 ;
      END
   END din0[10]
   PIN din0[11]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  143.04 0.0 143.42 0.38 ;
      END
   END din0[11]
   PIN din0[12]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  148.88 0.0 149.26 0.38 ;
      END
   END din0[12]
   PIN din0[13]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  154.72 0.0 155.1 0.38 ;
      END
   END din0[13]
   PIN din0[14]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  160.56 0.0 160.94 0.38 ;
      END
   END din0[14]
   PIN din0[15]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  166.4 0.0 166.78 0.38 ;
      END
   END din0[15]
   PIN din0[16]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  172.24 0.0 172.62 0.38 ;
      END
   END din0[16]
   PIN din0[17]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  178.08 0.0 178.46 0.38 ;
      END
   END din0[17]
   PIN din0[18]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  183.92 0.0 184.3 0.38 ;
      END
   END din0[18]
   PIN din0[19]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  189.76 0.0 190.14 0.38 ;
      END
   END din0[19]
   PIN din0[20]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  195.6 0.0 195.98 0.38 ;
      END
   END din0[20]
   PIN din0[21]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  201.44 0.0 201.82 0.38 ;
      END
   END din0[21]
   PIN din0[22]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  207.28 0.0 207.66 0.38 ;
      END
   END din0[22]
   PIN din0[23]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  213.12 0.0 213.5 0.38 ;
      END
   END din0[23]
   PIN din0[24]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  218.96 0.0 219.34 0.38 ;
      END
   END din0[24]
   PIN din0[25]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  224.8 0.0 225.18 0.38 ;
      END
   END din0[25]
   PIN din0[26]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  230.64 0.0 231.02 0.38 ;
      END
   END din0[26]
   PIN din0[27]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  236.48 0.0 236.86 0.38 ;
      END
   END din0[27]
   PIN din0[28]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  242.32 0.0 242.7 0.38 ;
      END
   END din0[28]
   PIN din0[29]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  248.16 0.0 248.54 0.38 ;
      END
   END din0[29]
   PIN din0[30]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  254.0 0.0 254.38 0.38 ;
      END
   END din0[30]
   PIN din0[31]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  259.84 0.0 260.22 0.38 ;
      END
   END din0[31]
   PIN din0[32]
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  265.68 0.0 266.06 0.38 ;
      END
   END din0[32]
   PIN addr0[0]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 124.53 0.38 124.91 ;
      END
   END addr0[0]
   PIN addr0[1]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 133.03 0.38 133.41 ;
      END
   END addr0[1]
   PIN addr0[2]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 138.67 0.38 139.05 ;
      END
   END addr0[2]
   PIN addr0[3]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 147.17 0.38 147.55 ;
      END
   END addr0[3]
   PIN addr0[4]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 153.075 0.38 153.455 ;
      END
   END addr0[4]
   PIN addr0[5]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 161.475 0.38 161.855 ;
      END
   END addr0[5]
   PIN addr0[6]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 166.95 0.38 167.33 ;
      END
   END addr0[6]
   PIN addr0[7]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 175.45 0.38 175.83 ;
      END
   END addr0[7]
   PIN addr0[8]
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 181.09 0.38 181.47 ;
      END
   END addr0[8]
   PIN csb0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 14.87 0.38 15.25 ;
      END
   END csb0
   PIN web0
      DIRECTION INPUT ;
      PORT
         LAYER met3 ;
         RECT  0.0 23.37 0.38 23.75 ;
      END
   END web0
   PIN clk0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  31.1 0.0 31.48 0.38 ;
      END
   END clk0
   PIN spare_wen0
      DIRECTION INPUT ;
      PORT
         LAYER met4 ;
         RECT  271.52 0.0 271.9 0.38 ;
      END
   END spare_wen0
   PIN dout0[0]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  143.79 0.0 144.17 0.38 ;
      END
   END dout0[0]
   PIN dout0[1]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  146.26 0.0 146.64 0.38 ;
      END
   END dout0[1]
   PIN dout0[2]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  149.57 0.0 149.95 0.38 ;
      END
   END dout0[2]
   PIN dout0[3]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  152.64 0.0 153.02 0.38 ;
      END
   END dout0[3]
   PIN dout0[4]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  155.41 0.0 155.79 0.38 ;
      END
   END dout0[4]
   PIN dout0[5]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  157.64 0.0 158.02 0.38 ;
      END
   END dout0[5]
   PIN dout0[6]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  158.755 0.0 159.135 0.38 ;
      END
   END dout0[6]
   PIN dout0[7]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  162.64 0.0 163.02 0.38 ;
      END
   END dout0[7]
   PIN dout0[8]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  163.79 0.0 164.17 0.38 ;
      END
   END dout0[8]
   PIN dout0[9]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  167.64 0.0 168.02 0.38 ;
      END
   END dout0[9]
   PIN dout0[10]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  168.79 0.0 169.17 0.38 ;
      END
   END dout0[10]
   PIN dout0[11]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  172.93 0.0 173.31 0.38 ;
      END
   END dout0[11]
   PIN dout0[12]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  173.79 0.0 174.17 0.38 ;
      END
   END dout0[12]
   PIN dout0[13]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  176.26 0.0 176.64 0.38 ;
      END
   END dout0[13]
   PIN dout0[14]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  178.79 0.0 179.17 0.38 ;
      END
   END dout0[14]
   PIN dout0[15]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  182.115 0.0 182.495 0.38 ;
      END
   END dout0[15]
   PIN dout0[16]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  184.61 0.0 184.99 0.38 ;
      END
   END dout0[16]
   PIN dout0[17]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  187.64 0.0 188.02 0.38 ;
      END
   END dout0[17]
   PIN dout0[18]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  190.45 0.0 190.83 0.38 ;
      END
   END dout0[18]
   PIN dout0[19]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  192.64 0.0 193.02 0.38 ;
      END
   END dout0[19]
   PIN dout0[20]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  193.79 0.0 194.17 0.38 ;
      END
   END dout0[20]
   PIN dout0[21]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  197.64 0.0 198.02 0.38 ;
      END
   END dout0[21]
   PIN dout0[22]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  198.79 0.0 199.17 0.38 ;
      END
   END dout0[22]
   PIN dout0[23]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  202.64 0.0 203.02 0.38 ;
      END
   END dout0[23]
   PIN dout0[24]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  203.79 0.0 204.17 0.38 ;
      END
   END dout0[24]
   PIN dout0[25]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  207.97 0.0 208.35 0.38 ;
      END
   END dout0[25]
   PIN dout0[26]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  208.79 0.0 209.17 0.38 ;
      END
   END dout0[26]
   PIN dout0[27]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  211.26 0.0 211.64 0.38 ;
      END
   END dout0[27]
   PIN dout0[28]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  213.85 0.0 214.23 0.38 ;
      END
   END dout0[28]
   PIN dout0[29]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  217.155 0.0 217.535 0.38 ;
      END
   END dout0[29]
   PIN dout0[30]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  220.17 0.0 220.55 0.38 ;
      END
   END dout0[30]
   PIN dout0[31]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  222.64 0.0 223.02 0.38 ;
      END
   END dout0[31]
   PIN dout0[32]
      DIRECTION OUTPUT ;
      PORT
         LAYER met4 ;
         RECT  226.335 0.0 226.715 0.38 ;
      END
   END dout0[32]
   PIN vccd1
      DIRECTION INOUT ;
      USE POWER ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met3 ;
         RECT  0.0 0.0 288.94 1.74 ;
         LAYER met4 ;
         RECT  0.0 0.0 1.74 502.86 ;
         LAYER met3 ;
         RECT  0.0 501.12 288.94 502.86 ;
         LAYER met4 ;
         RECT  287.2 0.0 288.94 502.86 ;
      END
   END vccd1
   PIN vssd1
      DIRECTION INOUT ;
      USE GROUND ; 
      SHAPE ABUTMENT ; 
      PORT
         LAYER met4 ;
         RECT  283.72 3.48 285.46 499.38 ;
         LAYER met3 ;
         RECT  3.48 3.48 285.46 5.22 ;
         LAYER met4 ;
         RECT  3.48 3.48 5.22 499.38 ;
         LAYER met3 ;
         RECT  3.48 497.64 285.46 499.38 ;
      END
   END vssd1
   OBS
   LAYER  met1 ;
      RECT  0.62 0.62 288.32 502.24 ;
   LAYER  met2 ;
      RECT  0.62 0.62 288.32 502.24 ;
   LAYER  met3 ;
      RECT  0.98 123.93 288.32 125.51 ;
      RECT  0.62 125.51 0.98 132.43 ;
      RECT  0.62 134.01 0.98 138.07 ;
      RECT  0.62 139.65 0.98 146.57 ;
      RECT  0.62 148.15 0.98 152.475 ;
      RECT  0.62 154.055 0.98 160.875 ;
      RECT  0.62 162.455 0.98 166.35 ;
      RECT  0.62 167.93 0.98 174.85 ;
      RECT  0.62 176.43 0.98 180.49 ;
      RECT  0.62 15.85 0.98 22.77 ;
      RECT  0.62 24.35 0.98 123.93 ;
      RECT  0.62 2.34 0.98 14.27 ;
      RECT  0.62 182.07 0.98 500.52 ;
      RECT  0.98 2.34 2.88 2.88 ;
      RECT  0.98 2.88 2.88 5.82 ;
      RECT  0.98 5.82 2.88 123.93 ;
      RECT  2.88 2.34 286.06 2.88 ;
      RECT  2.88 5.82 286.06 123.93 ;
      RECT  286.06 2.34 288.32 2.88 ;
      RECT  286.06 2.88 288.32 5.82 ;
      RECT  286.06 5.82 288.32 123.93 ;
      RECT  0.98 125.51 2.88 497.04 ;
      RECT  0.98 497.04 2.88 499.98 ;
      RECT  0.98 499.98 2.88 500.52 ;
      RECT  2.88 125.51 286.06 497.04 ;
      RECT  2.88 499.98 286.06 500.52 ;
      RECT  286.06 125.51 288.32 497.04 ;
      RECT  286.06 497.04 288.32 499.98 ;
      RECT  286.06 499.98 288.32 500.52 ;
   LAYER  met4 ;
      RECT  78.2 0.98 79.78 502.24 ;
      RECT  79.78 0.62 84.04 0.98 ;
      RECT  85.62 0.62 89.88 0.98 ;
      RECT  91.46 0.62 95.72 0.98 ;
      RECT  97.3 0.62 101.56 0.98 ;
      RECT  103.14 0.62 107.4 0.98 ;
      RECT  108.98 0.62 113.24 0.98 ;
      RECT  114.82 0.62 119.08 0.98 ;
      RECT  120.66 0.62 124.92 0.98 ;
      RECT  126.5 0.62 130.76 0.98 ;
      RECT  132.34 0.62 136.6 0.98 ;
      RECT  138.18 0.62 142.44 0.98 ;
      RECT  231.62 0.62 235.88 0.98 ;
      RECT  237.46 0.62 241.72 0.98 ;
      RECT  243.3 0.62 247.56 0.98 ;
      RECT  249.14 0.62 253.4 0.98 ;
      RECT  254.98 0.62 259.24 0.98 ;
      RECT  260.82 0.62 265.08 0.98 ;
      RECT  32.08 0.62 78.2 0.98 ;
      RECT  266.66 0.62 270.92 0.98 ;
      RECT  144.77 0.62 145.66 0.98 ;
      RECT  147.24 0.62 148.28 0.98 ;
      RECT  150.55 0.62 152.04 0.98 ;
      RECT  153.62 0.62 154.12 0.98 ;
      RECT  156.39 0.62 157.04 0.98 ;
      RECT  159.735 0.62 159.96 0.98 ;
      RECT  161.54 0.62 162.04 0.98 ;
      RECT  164.77 0.62 165.8 0.98 ;
      RECT  169.77 0.62 171.64 0.98 ;
      RECT  174.77 0.62 175.66 0.98 ;
      RECT  177.24 0.62 177.48 0.98 ;
      RECT  179.77 0.62 181.515 0.98 ;
      RECT  183.095 0.62 183.32 0.98 ;
      RECT  185.59 0.62 187.04 0.98 ;
      RECT  188.62 0.62 189.16 0.98 ;
      RECT  191.43 0.62 192.04 0.98 ;
      RECT  194.77 0.62 195.0 0.98 ;
      RECT  196.58 0.62 197.04 0.98 ;
      RECT  199.77 0.62 200.84 0.98 ;
      RECT  204.77 0.62 206.68 0.98 ;
      RECT  209.77 0.62 210.66 0.98 ;
      RECT  212.24 0.62 212.52 0.98 ;
      RECT  214.83 0.62 216.555 0.98 ;
      RECT  218.135 0.62 218.36 0.98 ;
      RECT  221.15 0.62 222.04 0.98 ;
      RECT  223.62 0.62 224.2 0.98 ;
      RECT  227.315 0.62 230.04 0.98 ;
      RECT  2.34 0.62 30.5 0.98 ;
      RECT  272.5 0.62 286.6 0.98 ;
      RECT  79.78 0.98 283.12 2.88 ;
      RECT  79.78 2.88 283.12 499.98 ;
      RECT  79.78 499.98 283.12 502.24 ;
      RECT  283.12 0.98 286.06 2.88 ;
      RECT  283.12 499.98 286.06 502.24 ;
      RECT  286.06 0.98 286.6 2.88 ;
      RECT  286.06 2.88 286.6 499.98 ;
      RECT  286.06 499.98 286.6 502.24 ;
      RECT  2.34 0.98 2.88 2.88 ;
      RECT  2.34 2.88 2.88 499.98 ;
      RECT  2.34 499.98 2.88 502.24 ;
      RECT  2.88 0.98 5.82 2.88 ;
      RECT  2.88 499.98 5.82 502.24 ;
      RECT  5.82 0.98 78.2 2.88 ;
      RECT  5.82 2.88 78.2 499.98 ;
      RECT  5.82 499.98 78.2 502.24 ;
   END
END    sram_32b_256_1rw_sky130
END    LIBRARY
